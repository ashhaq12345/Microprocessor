CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
48 C:\Program Files\CircuitMaker 2000 Trial\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
28
13 Logic Switch~
5 164 338 0 1 11
0 41
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5305 0 0
2
41840 0
0
13 Logic Switch~
5 211 340 0 10 11
0 42 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
34 0 0
2
41840 0
0
13 Logic Switch~
5 259 338 0 1 11
0 43
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
969 0 0
2
41840 0
0
13 Logic Switch~
5 303 337 0 10 11
0 44 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8402 0 0
2
41840 0
0
13 Logic Switch~
5 39 102 0 10 11
0 45 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3751 0 0
2
5.8967e-315 0
0
13 Logic Switch~
5 61 186 0 10 11
0 47 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4292 0 0
2
5.8967e-315 0
0
14 Logic Display~
6 621 982 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6118 0 0
2
41840.1 0
0
14 Logic Display~
6 653 983 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
34 0 0
2
41840.1 0
0
14 Logic Display~
6 681 984 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6357 0 0
2
41840.1 0
0
14 Logic Display~
6 712 988 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
319 0 0
2
41840.1 0
0
7 74LS173
129 259 687 0 14 29
0 15 6 6 16 17 18 19 20 5
5 11 12 13 14
0
0 0 4848 782
6 74F173
-21 -51 21 -43
2 U9
48 -2 62 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
3976 0 0
2
41840.1 0
0
6 PROM32
80 756 169 0 14 29
0 15 30 29 28 27 26 25 24 23
22 21 4 2 3
0
0 0 4848 0
6 PROM32
-21 -19 21 -11
3 U11
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 4 5 6 7 9 10
11 12 13 14 15 1 2 3 4 5
6 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
7634 0 0
2
41840 0
0
PPPPPPPPPNPOCKAAAAAAAAAAAAAAAAAAAPAPPPAAAAAAAAAAAAAAAAAAAAAAAAAA
14 Logic Display~
6 27 363 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
523 0 0
2
41840 0
0
14 Logic Display~
6 55 364 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6748 0 0
2
41840 0
0
14 Logic Display~
6 86 365 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6901 0 0
2
41840 0
0
14 Logic Display~
6 122 364 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
842 0 0
2
41840 0
0
7 74LS173
129 655 794 0 14 29
0 15 2 2 16 17 18 19 20 3
3 31 32 33 34
0
0 0 4848 782
6 74F173
-21 -51 21 -43
3 U10
45 -2 66 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
3277 0 0
2
41840 0
0
7 74LS173
129 626 655 0 14 29
0 15 36 36 16 17 18 19 20 35
35 17 18 19 20
0
0 0 4848 782
6 74F173
-21 -51 21 -43
2 U8
48 -2 62 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
4212 0 0
2
41840 0
0
7 74LS173
129 253 464 0 14 29
0 15 40 40 16 41 42 43 44 39
39 17 18 19 20
0
0 0 4848 782
6 74F173
-21 -51 21 -43
2 U5
48 -2 62 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
4720 0 0
2
41840 0
0
7 74LS181
132 701 894 0 22 45
0 25 24 23 22 17 18 19 20 31
32 33 34 21 4 49 50 51 52 7
8 9 10
0
0 0 4848 270
6 74F181
-21 -69 21 -61
2 U7
66 -2 80 6
0
16 DVCC=24;DGND=12;
192 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 3 4 5 6 19 21 23 2 18
20 22 1 7 8 16 14 17 15 13
11 10 9 3 4 5 6 19 21 23
2 18 20 22 1 7 8 16 14 17
15 13 11 10 9 0
65 0 0 512 1 0 0 0
1 U
5551 0 0
2
5.8967e-315 0
0
7 74LS173
129 691 465 0 14 29
0 15 38 38 16 17 18 19 20 37
37 17 18 19 20
0
0 0 4848 782
6 74F173
-21 -51 21 -43
2 U6
48 -2 62 6
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
6986 0 0
2
5.8967e-315 0
0
6 PROM32
80 532 172 0 14 29
0 15 30 29 28 27 26 40 39 38
37 36 35 6 5
0
0 0 4848 0
6 PROM32
-21 -19 21 -11
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 4 5 6 7 9 10
11 12 13 14 15 1 2 3 4 5
6 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
8745 0 0
2
5.8967e-315 0
0
DPJPPPDPLPOPOPPOAAAAAAAAAAAAAAAAAPAPPPAAAAAAAAAAAAAAAAAAAAAAAAAA
6 74LS93
109 411 77 0 8 17
0 15 15 29 53 54 55 56 30
0
0 0 4848 0
6 74LS93
-21 -35 21 -27
2 U3
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 512 1 0 0 0
1 U
9592 0 0
2
5.8967e-315 0
0
14 NO PushButton~
191 105 97 0 2 5
0 46 45
0
0 0 4720 0
0
2 S2
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
8748 0 0
2
5.8967e-315 5.30499e-315
0
9 2-In AND~
219 190 113 0 3 22
0 45 46 15
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
7168 0 0
2
5.8967e-315 5.26354e-315
0
9 2-In AND~
219 212 197 0 3 22
0 47 48 16
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
631 0 0
2
5.8967e-315 0
0
14 NO PushButton~
191 127 181 0 2 5
0 48 47
0
0 0 4720 0
0
2 S1
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
9466 0 0
2
5.8967e-315 0
0
6 74LS93
109 324 169 0 8 17
0 15 15 16 26 29 28 27 26
0
0 0 4848 0
6 74LS93
-21 -35 21 -27
2 U1
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
3266 0 0
2
5.8967e-315 0
0
126
3 13 2 0 0 12416 0 17 12 0 0 5
644 758
644 699
796 699
796 196
788 196
14 0 3 0 0 8192 0 12 0 0 24 4
788 205
861 205
861 397
866 397
12 0 4 0 0 8192 0 12 0 0 22 4
788 187
889 187
889 415
894 415
10 14 5 0 0 12416 0 11 22 0 0 5
239 727
239 751
577 751
577 208
564 208
3 13 6 0 0 8320 0 11 22 0 0 5
248 651
248 533
587 533
587 199
564 199
9 10 5 0 0 0 0 11 11 0 0 3
230 727
230 727
239 727
19 1 7 0 0 8320 0 20 7 0 0 6
676 934
676 957
608 957
608 1008
621 1008
621 1000
20 1 8 0 0 4224 0 20 8 0 0 4
667 934
667 1009
653 1009
653 1001
21 1 9 0 0 12416 0 20 9 0 0 6
658 934
658 964
668 964
668 1010
681 1010
681 1002
22 1 10 0 0 8320 0 20 10 0 0 6
649 934
649 968
699 968
699 1014
712 1014
712 1006
11 1 11 0 0 12416 0 11 13 0 0 4
266 721
266 746
27 746
27 381
12 1 12 0 0 12416 0 11 14 0 0 4
275 721
275 741
55 741
55 382
13 1 13 0 0 12416 0 11 15 0 0 4
284 721
284 736
86 736
86 383
14 1 14 0 0 12416 0 11 16 0 0 4
293 721
293 731
122 731
122 382
2 3 6 0 0 0 0 11 11 0 0 3
239 651
239 651
248 651
1 3 15 0 0 20480 0 11 25 0 0 7
230 657
230 513
199 513
199 365
243 365
243 113
211 113
4 3 16 0 0 20480 0 11 26 0 0 7
257 657
257 508
204 508
204 360
241 360
241 197
233 197
5 0 17 0 0 8192 0 11 0 0 107 5
266 657
266 632
370 632
370 658
375 658
6 0 18 0 0 8192 0 11 0 0 106 5
275 657
275 637
422 637
422 662
427 662
7 0 19 0 0 8192 0 11 0 0 105 5
284 657
284 642
474 642
474 661
479 661
8 0 20 0 0 8192 0 11 0 0 104 3
293 657
293 647
527 647
14 0 4 0 0 12416 0 20 0 0 0 5
739 928
739 938
894 938
894 400
899 400
0 10 3 0 0 4224 0 0 17 24 0 9
866 403
640 403
640 615
675 615
675 724
606 724
606 842
635 842
635 834
0 0 3 0 0 0 0 0 0 0 0 2
866 389
866 407
0 13 21 0 0 8320 0 0 20 30 0 5
942 433
768 433
768 942
748 942
748 928
4 0 22 0 0 4224 0 20 0 0 31 5
721 864
721 514
960 514
960 425
965 425
3 0 23 0 0 4224 0 20 0 0 32 5
730 864
730 509
980 509
980 433
985 433
2 0 24 0 0 4224 0 20 0 0 36 3
739 864
739 447
1006 447
1 0 25 0 0 4224 0 20 0 0 35 3
748 864
748 455
1025 455
11 0 21 0 0 0 0 12 0 0 39 4
788 178
942 178
942 442
947 442
10 0 22 0 0 0 0 12 0 0 38 4
788 169
965 169
965 442
970 442
9 0 23 0 0 0 0 12 0 0 37 4
788 160
985 160
985 439
990 439
8 0 24 0 0 0 0 12 0 0 36 4
788 151
1001 151
1001 440
1006 440
7 0 25 0 0 0 0 12 0 0 35 4
788 142
1020 142
1020 440
1025 440
0 0 25 0 0 0 0 0 0 0 0 2
1025 436
1025 460
0 0 24 0 0 0 0 0 0 0 0 2
1006 437
1006 458
0 0 23 0 0 0 0 0 0 0 0 2
990 435
990 456
0 0 22 0 0 0 0 0 0 0 0 2
970 435
970 454
0 0 21 0 0 0 0 0 0 0 0 2
947 433
947 454
9 10 3 0 0 0 0 17 17 0 0 3
626 834
626 834
635 834
2 3 2 0 0 0 0 17 17 0 0 3
635 758
635 758
644 758
4 4 16 0 0 0 0 17 18 0 0 6
653 764
653 704
567 704
567 611
624 611
624 625
1 1 15 0 0 0 0 18 17 0 0 6
597 625
597 615
572 615
572 735
626 735
626 764
6 6 26 0 0 12416 0 22 12 0 0 6
500 208
485 208
485 248
695 248
695 205
724 205
5 5 27 0 0 12416 0 22 12 0 0 6
500 199
475 199
475 243
700 243
700 196
724 196
4 4 28 0 0 12416 0 22 12 0 0 6
500 190
470 190
470 238
705 238
705 187
724 187
3 3 29 0 0 12416 0 22 12 0 0 6
500 181
490 181
490 233
710 233
710 178
724 178
2 2 30 0 0 12416 0 22 12 0 0 6
500 172
470 172
470 101
705 101
705 169
724 169
1 1 15 0 0 0 0 22 12 0 0 6
494 136
490 136
490 111
710 111
710 133
718 133
11 5 17 0 0 4096 0 21 20 0 0 4
698 499
698 754
712 754
712 858
12 6 18 0 0 4096 0 21 20 0 0 4
707 499
707 840
703 840
703 858
13 7 19 0 0 4096 0 21 20 0 0 4
716 499
716 850
694 850
694 858
14 8 20 0 0 4096 0 21 20 0 0 4
725 499
725 845
685 845
685 858
11 9 31 0 0 12416 0 17 20 0 0 4
662 828
662 840
676 840
676 858
12 10 32 0 0 12416 0 17 20 0 0 4
671 828
671 840
667 840
667 858
13 11 33 0 0 8320 0 17 20 0 0 4
680 828
680 845
658 845
658 858
14 12 34 0 0 8320 0 17 20 0 0 4
689 828
689 850
649 850
649 858
5 0 17 0 0 8192 0 17 0 0 107 3
662 764
662 741
375 741
6 0 18 0 0 0 0 17 0 0 106 3
671 764
671 744
427 744
7 0 19 0 0 0 0 17 0 0 105 3
680 764
680 748
479 748
8 0 20 0 0 0 0 17 0 0 104 3
689 764
689 754
527 754
9 12 35 0 0 12416 0 18 22 0 0 5
597 695
597 699
577 699
577 190
564 190
2 11 36 0 0 4224 0 18 22 0 0 3
606 619
606 181
564 181
9 10 37 0 0 12416 0 21 22 0 0 5
662 505
662 509
582 509
582 172
564 172
2 9 38 0 0 4224 0 21 22 0 0 3
671 429
671 163
564 163
9 8 39 0 0 12416 0 19 22 0 0 5
224 504
224 518
577 518
577 154
564 154
2 7 40 0 0 8320 0 19 22 0 0 5
233 428
233 228
572 228
572 145
564 145
2 3 36 0 0 128 0 18 18 0 0 2
606 619
615 619
10 9 35 0 0 128 0 18 18 0 0 2
606 695
597 695
4 0 16 0 0 8320 0 18 0 0 123 6
624 625
624 389
239 389
239 202
253 202
253 197
1 0 15 0 0 4224 0 18 0 0 118 4
597 625
597 116
220 116
220 113
11 0 17 0 0 0 0 18 0 0 107 3
633 689
633 729
375 729
12 0 18 0 0 0 0 18 0 0 106 3
642 689
642 707
427 707
13 0 19 0 0 0 0 18 0 0 105 3
651 689
651 713
479 713
14 0 20 0 0 0 0 18 0 0 104 3
660 689
660 717
527 717
5 0 17 0 0 0 0 18 0 0 107 3
633 625
633 590
375 590
6 0 18 0 0 0 0 18 0 0 106 3
642 625
642 592
427 592
7 0 19 0 0 0 0 18 0 0 105 3
651 625
651 596
479 596
8 0 20 0 0 0 0 18 0 0 104 3
660 625
660 599
527 599
1 0 15 0 0 0 0 21 0 0 118 4
662 435
662 108
227 108
227 113
11 0 17 0 0 8192 0 21 0 0 107 3
698 499
698 561
375 561
12 0 18 0 0 0 0 21 0 0 106 3
707 499
707 565
427 565
13 0 19 0 0 0 0 21 0 0 105 3
716 499
716 570
479 570
14 0 20 0 0 0 0 21 0 0 104 3
725 499
725 573
527 573
10 9 37 0 0 0 0 21 21 0 0 2
671 505
662 505
3 2 38 0 0 0 0 21 21 0 0 2
680 429
671 429
4 0 16 0 0 0 0 21 0 0 123 6
689 435
689 202
568 202
568 223
262 223
262 197
5 0 17 0 0 0 0 21 0 0 107 3
698 435
698 421
375 421
6 0 18 0 0 0 0 21 0 0 106 3
707 435
707 418
427 418
7 0 19 0 0 0 0 21 0 0 105 3
716 435
716 413
479 413
8 0 20 0 0 0 0 21 0 0 104 3
725 435
725 410
527 410
1 0 15 0 0 0 0 19 0 0 118 4
224 434
224 355
238 355
238 113
11 0 17 0 0 0 0 19 0 0 107 3
260 498
260 529
375 529
12 0 18 0 0 0 0 19 0 0 106 3
269 498
269 522
427 522
13 0 19 0 0 0 0 19 0 0 105 3
278 498
278 514
479 514
14 0 20 0 0 0 0 19 0 0 104 3
287 498
287 508
527 508
9 10 39 0 0 0 0 19 19 0 0 2
224 504
233 504
2 3 40 0 0 0 0 19 19 0 0 2
233 428
242 428
4 0 16 0 0 0 0 19 0 0 123 4
251 434
251 358
244 358
244 197
5 1 41 0 0 4224 0 19 1 0 0 5
260 434
260 351
185 351
185 338
176 338
6 1 42 0 0 4224 0 19 2 0 0 5
269 434
269 348
232 348
232 340
223 340
7 1 43 0 0 4224 0 19 3 0 0 3
278 434
278 338
271 338
8 1 44 0 0 4224 0 19 4 0 0 5
287 434
287 348
324 348
324 337
315 337
0 0 20 0 0 4224 0 0 0 0 0 2
527 284
527 935
0 0 19 0 0 4224 0 0 0 0 0 2
479 281
479 936
0 0 18 0 0 4224 0 0 0 0 0 2
427 280
427 937
0 0 17 0 0 4224 0 0 0 0 0 2
375 278
375 936
0 1 15 0 0 0 0 0 22 118 0 3
265 113
265 136
494 136
8 6 26 0 0 128 0 28 22 0 0 4
356 187
481 187
481 208
500 208
7 5 27 0 0 128 0 28 22 0 0 4
356 178
486 178
486 199
500 199
6 4 28 0 0 128 0 28 22 0 0 4
356 169
476 169
476 190
500 190
5 3 29 0 0 128 0 28 22 0 0 4
356 160
481 160
481 181
500 181
8 2 30 0 0 128 0 23 22 0 0 4
443 95
486 95
486 172
500 172
5 3 29 0 0 0 0 28 23 0 0 4
356 160
365 160
365 86
373 86
2 0 15 0 0 0 0 23 0 0 118 3
379 77
251 77
251 113
0 1 15 0 0 0 0 0 23 118 0 3
236 113
236 68
379 68
4 8 26 0 0 0 0 28 28 0 0 6
286 187
282 187
282 202
364 202
364 187
356 187
3 2 15 0 0 0 0 25 28 0 0 4
211 113
273 113
273 169
292 169
3 1 15 0 0 0 0 25 28 0 0 4
211 113
278 113
278 160
292 160
2 1 45 0 0 4096 0 24 5 0 0 4
88 105
60 105
60 102
51 102
1 1 45 0 0 12416 0 5 25 0 0 6
51 102
84 102
84 113
153 113
153 104
166 104
1 2 46 0 0 4224 0 24 25 0 0 4
122 105
158 105
158 122
166 122
3 3 16 0 0 0 0 26 28 0 0 4
233 197
273 197
273 178
286 178
2 1 47 0 0 4096 0 27 6 0 0 4
110 189
82 189
82 186
73 186
1 1 47 0 0 12416 0 6 26 0 0 6
73 186
106 186
106 197
175 197
175 188
188 188
1 2 48 0 0 4224 0 27 26 0 0 4
144 189
180 189
180 206
188 206
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
810 881 855 905
820 889 844 905
3 ALU
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
741 784 794 808
751 792 783 808
4 Temp
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
701 645 730 669
711 653 719 669
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
765 453 794 477
775 461 783 477
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
156 458 217 482
166 466 206 482
5 Input
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-06 1e-07 1e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
